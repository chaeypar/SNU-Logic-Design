`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:39:56 05/18/2023 
// Design Name: 
// Module Name:    gated_RS_latch 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gated_RS_latch(
    input R,
    input S,
    input E,
    output Q,
    output Qinv
    );
	
	reg r, s;
	
	always @(E or R or S)
		begin
			r = R & E;
			s = S & E;
		end
	RS_latch T1(.R(r), .S(s), .Q(Q), .Qinv(Qinv));
	
endmodule

























































































































































































































































































































































































































































































































































































































































